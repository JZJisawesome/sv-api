module hello();
    wire b;
endmodule

module top();
    wire a;
    hello h();
endmodule
