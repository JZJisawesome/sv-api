/*
 * File:    TODO.sv
 * Brief:   TODO
 *
 * Copyright (C) TODO John Jekel
 * See the LICENSE file at the root of the project for licensing info.
 *
 * TODO longer description
 *
*/

module hello();
    wire b;
endmodule

module top();
    reg a;
    hello h();
endmodule
