module hello();
    wire b;
endmodule

module top();
    reg a;
    hello h();
endmodule
